//
// eJ32 - Java Forth Machine - Load/Store Unit
//
`include "../source/eJ32_if.sv"

module EJ32_LS #(
    parameter TIB      = 'h1000,          ///> input buffer address
    parameter OBUF     = 'h1400,          ///> output buffer address
    parameter DSZ      = 32,              ///> 32-bit data width
    parameter ASZ      = 17               ///> 128K address space
    ) (
    EJ32_CTL ctl,
    input  `U1 ls_en,
    input  `U8 data,                      ///> data from memory bus
    input  `DU s,                         ///> NOS
    output `U1 ls_asel_o,
    output `IU ls_addr_o,                 ///> address to memory bus
    output `U8 data_o,                    ///> data to memory bus
    output `U1 dwe_o                      ///> data write enable
    );
    import ej32_pkg::*;
    /// @defgroup Registers
    /// @{
    // instruction
    `IU  a;                     ///> memory address
    `IU  asel;
    // IO
    `U2  dsel;                  ///> 32-bit, 4-to-1 mux, byte select
    `IU  ibuf, obuf;            ///> input, output buffer pointers
    /// @}
    /// @defgroup Next Register
    /// @{
    `DU t_n;                    ///> TOS
    `IU a_n;                    ///> data address
    `IU asel_n;                 ///> address select
    `U8 data_n;
    `U2 dsel_n;                 ///> 32-bit, 4-to-1 mux, byte select
    /// @}
    /// @defgroup Wires
    /// @{
    // instruction
    opcode_t code;              ///> shadow ctl.code
    `U3  phase;                 ///> FSM phase (aka state)
    `U1 a_x;                    ///> address controls
    `IU a_d;                    ///> 2-byte merged address
    // data stack
    `DU t;                      ///> shadow TOS
    `U1 t_x;
    `DU t_d;                    ///> 4-byte merged data
    // memory & IO buffers
    `U8 d8x4[4];                ///> 4-to-1 byte select
    `U1 dwe, dsel_x;            ///> data/addr bus controls
    `U1 ibuf_x, obuf_x;         ///> input/output buffer controls
    /// @}

    task TOS(input `DU v);  t_n = v; `SET(t_x);   endtask;   ///> update TOS
    task SETA(input `IU a); a_n = a; `SET(a_x);   endtask;   ///> build addr ptr
    task MEM(input `IU a); SETA(a); `SET(asel_n); endtask;   ///> fetch from memory, data returns next cycle
    task DW(input `U3 n); dsel_n = n; `SET(dwe); `SET(dsel_x); endtask;   ///> data write n-th byte
    ///
    /// wires to reduce verbosity
    ///
    assign code     = ctl.code;               ///> input from ej32 control
    assign phase    = ctl.phase;
    assign t        = ctl.t;
    assign ls_addr_o= a;                      ///> memory address
    assign ls_asel_o= asel;
    assign data_o   = data_n;                 ///> data sent to memory bus
    assign dwe_o    = dwe;                    ///> data write enable
    assign d8x4     =                         ///> 4-to-1 Big-Endian
        {t[31:24],t[23:16],t[15:8],t[7:0]};
    assign data_n   = d8x4[dsel];             ///> data byte select (Big-Endian)
    ///
    /// wires to external modules
    ///
    assign a_d    = {a[ASZ-9:0], data};       ///> merge lowest byte into addr
    assign t_d    = {t[DSZ-9:0], data};       ///> merge lowest byte into TOS
    ///
    /// combinational
    ///
    task INIT();
        t_n       = {DSZ{1'b0}};  /// TOS
        t_x       = 1'b0;
        a_n       = {ASZ{1'b0}};  /// default to clear address
        a_x       = 1'b0;
        asel_n    = 1'b0;         /// address default to program counter
        dsel_x    = 1'b0;         /// data bus
        dsel_n    = 3;
        dwe       = 1'b0;         /// data write
        ibuf_x    = 1'b0;
        obuf_x    = 1'b0;
    endtask: INIT

    always_comb begin
        INIT();
        case (code)
        iaload:
            case (phase)
            0: MEM(`XDA(t));
            1: begin MEM(a + 1); TOS(`X8D(data)); end
            2: begin MEM(a + 1); TOS(t_d); end
            3: begin MEM(a + 1); TOS(t_d); end
            4: TOS(t_d);
            endcase
        baload:
            case (phase)
            0: MEM(`XDA(t));
            1: TOS(`X8D(data));
            endcase
        saload:
            case (phase)
            0: MEM(`XDA(t));
            1: begin MEM(a + 1); TOS(`X8D(data)); end
            2: TOS(t_d);
            endcase
        iastore:
            case (phase)
            0: begin MEM(`XDA(s)); `SET(dsel_x); dsel_n = 0; end
            1: begin MEM(a + 1); DW(1); end
            2: begin MEM(a + 1); DW(2); end
            3: begin MEM(a + 1); DW(3); end
            4: DW(3);                          // CC: reset a?
            endcase
        bastore:
            case (phase)
            0: MEM(`XDA(s));
            1: DW(3);                          // CC: reset a?
            endcase
        sastore:
            case (phase)                       // CC: logic changed from Dr. Ting's
            0: begin MEM(`XDA(s)); `SET(dsel_x); dsel_n = 2; end
            1: begin MEM(a + 1); DW(3); end
            2: DW(3);
            endcase
        iinc:
            case (phase)                       // CC: logic changed from Dr. Ting's
            0: MEM(`XDA(s));
            1: `SET(asel_n);
            2: begin TOS(s); DW(0); end
            endcase
        ldi: 
            case (phase)
            1: TOS(t_d);
            2: TOS(t_d);
            3: TOS(t_d);
            endcase
        get:
            case (phase)
            0: MEM(ibuf);
            1: begin TOS(`X8D(data)); `SET(ibuf_x); end
            endcase
        put:
            case (phase)
            0: begin MEM(obuf); `SET(dsel_x); end
            1: begin DW(3);     `SET(obuf_x); end
            endcase
        endcase
    end // always_comb

    always_ff @(posedge ctl.clk, posedge ctl.rst) begin
        if (ctl.rst) begin
            asel  <= 1'b0;
            dsel  <= 3;
            ibuf  <= TIB;
            obuf  <= OBUF;
            a     <= {ASZ{1'b0}};
        end
        else if (ctl.clk && ls_en) begin
            asel <= asel_n;
            if (t_x)     ctl.t    <= t_n;
            if (a_x)     a        <= a_n;
            if (dsel_x)  dsel     <= dsel_n;
            if (ibuf_x)  ibuf     <= ibuf + 1;
            if (obuf_x)  obuf     <= obuf + 1;
        end
    end // always_ff @ (posedge clk, posedge rst)
endmodule: EJ32_LS
